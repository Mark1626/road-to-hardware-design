module thruwire(
  input  wire i_in,
  output wire o_out
);

  assign o_out = i_in;

endmodule
